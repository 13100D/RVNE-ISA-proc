module rvne(input [31:0] instruction);
    wire [31:0] [31:0] regFile;
    
endmodule